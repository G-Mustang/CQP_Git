// ss1 testbench code
