// ss1 rtl code
//

module ss1;

initial begin
    $display("ff");
    $display("f1");
    $display("f2");
    $display("f3");
    $display("f4");
end

endmodule
