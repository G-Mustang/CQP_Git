// ss2 testbench code
