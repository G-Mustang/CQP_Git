// ss1 rtl code
//

module ss1;

initial begin
    $display("ff");
end

endmodule
