// ss1 rtl code
//

module ss1;

initial begin

end

endmodule
