// ss3 testbench code
