// ss2 rtl code
//
module ss2;

initial begin
    $display("aaaa");
end

endmodule
