// ss3 rtl code
//

module ss3;

initial begin
    $display("fff");
end

endmodule
